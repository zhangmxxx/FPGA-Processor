module bcd7seg(input [7:0] b, output reg [7:0] h);
  always @(*) begin
    case(b)
      8'd0: h = 8'b11000000; 
      8'd1: h = 8'b11111001; 
      8'd2: h = 8'b10100100; 
      8'd3: h = 8'b10110000; 
      8'd4: h = 8'b10011001; 
      8'd5: h = 8'b10010010; 
      8'd6: h = 8'b10000010; 
      8'd7: h = 8'b11111000; 
      8'd8: h = 8'b10000000;
      8'd9: h = 8'b10010000;
      8'd10: h = 8'b10001000;
      8'd11: h = 8'b10000011;
      8'd12: h = 8'b11000110;     
      8'd13: h = 8'b10100001;  
      8'd14: h = 8'b10000110;
      8'd15: h = 8'b10001110;
      default: h = 8'b11111111;
    endcase
  end  
endmodule